// Auto-assembled from src .sv files by copy_src_sv_to_fpga_sv.sh

// =======================
// The Tiny Tapeout module
// =======================

module tt_um_template (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
       // The FPGA is based on TinyTapeout 3 which has no bidirectional I/Os (vs. TT6 for the ASIC).
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

   // Parameters for Memory Sizing and UART Baud
   localparam int unsigned COUNTER_WIDTH = 24;       // Width of the clock counters in the UART RX and TX modules
   localparam int unsigned IMEM_BYTE_ADDR_WIDTH = 6; // 64 bytes / 16 words of I-Memory
   localparam int unsigned DMEM_BYTE_ADDR_WIDTH = 4; // 16 bytes /  4 words of D-Memory

   // CPU Reset
   wire reset;

   // User Interface
   wire rst = ! rst_n | ui_in[7]; // Provide a dedicated button input for RESET
   wire rx_in = ui_in[2];         // Should be wired to Pin 2 of the USBUART Pmod (data from host to Pmod)
   wire tx_out;
   assign uo_out[7] = rst;        // Feedback of RST button, intended to use with LED
   assign uo_out[6] = reset;      // Feedback of CPU reset, indicates if UART controller is in write mode (reset = 1) or read mode (reset = 0)
   assign uo_out[5] = ~rx_in;     // Feedback of RX line, intended to use with LED
   assign uo_out[4] = ~tx_out;    // Feedback of TX line, intended to use with LED
   assign uo_out[3] = 1'b0;       // Unused
   assign uo_out[2] = tx_out;     // Should be wired to Pin 3 of the USBUART Pmod (data from Pmod to host)
   assign uo_out[1] = 1'b0;       // Unused
   assign uo_out[0] = 1'b0;       // Unused

   // I-Memory Interface
   logic imem_rd_en;
   logic [IMEM_BYTE_ADDR_WIDTH-3:0] imem_rd_addr;
   logic [31:0] imem_rd_data;

   // D-Memory Interface
   logic dmem_rd_en, dmem_wr_en;
   logic [DMEM_BYTE_ADDR_WIDTH-3:0] dmem_addr;
   logic [3:0] dmem_wr_byte_en;
   logic [31:0] dmem_wr_data, dmem_rd_data;

   // UART Module
   uart_top #(
      .COUNTER_WIDTH(COUNTER_WIDTH),
      .IMEM_BYTE_ADDR_WIDTH(IMEM_BYTE_ADDR_WIDTH),
      .DMEM_BYTE_ADDR_WIDTH(DMEM_BYTE_ADDR_WIDTH))
   uart_top0 (
      .clk(clk),
      .rst(rst),
      .rx_in(rx_in),
      .tx_out(tx_out),
      .cpu_rst(reset),
      .imem_rd_en(imem_rd_en),
      .imem_rd_addr(imem_rd_addr),
      .imem_rd_data(imem_rd_data),
      .dmem_rd_en(dmem_rd_en),
      .dmem_wr_en(dmem_wr_en),
      .dmem_addr(dmem_addr),
      .dmem_wr_byte_en(dmem_wr_byte_en),
      .dmem_wr_data(dmem_wr_data),
      .dmem_rd_data(dmem_rd_data));

// ---------- Generated Code Inlined Here (before 1st \TLV) ----------
// Generated by SandPiper(TM) 1.14-2022/10/10-beta-Pro from Redwood EDA, LLC.
// (Installed here: /usr/local/mono/sandpiper/distro.)
// Redwood EDA, LLC does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


// For silencing unused signal messages.
`define BOGUS_USE(ignore)


genvar digit, input_label, leds, switch, xreg;


//
// Signals declared top-level.
//

// For $slideswitch.
logic [7:0] L0_slideswitch_a0;

// For $sseg_decimal_point_n.
logic L0_sseg_decimal_point_n_a0;

// For $sseg_digit_n.
logic [7:0] L0_sseg_digit_n_a0;

// For $sseg_segment_n.
logic [6:0] L0_sseg_segment_n_a0;

// For /fpga_pins/fpga|cpu$alu_op1.
logic [31:0] FpgaPins_Fpga_CPU_alu_op1_a2,
             FpgaPins_Fpga_CPU_alu_op1_a3;

// For /fpga_pins/fpga|cpu$alu_op2.
logic [31:0] FpgaPins_Fpga_CPU_alu_op2_a2,
             FpgaPins_Fpga_CPU_alu_op2_a3;

// For /fpga_pins/fpga|cpu$funct3.
logic [2:0] FpgaPins_Fpga_CPU_funct3_a1;

// For /fpga_pins/fpga|cpu$funct7.
logic [6:0] FpgaPins_Fpga_CPU_funct7_a1;

// For /fpga_pins/fpga|cpu$imm.
logic [31:0] FpgaPins_Fpga_CPU_imm_a1,
             FpgaPins_Fpga_CPU_imm_a2;

// For /fpga_pins/fpga|cpu$inc_pc.
logic [31:0] FpgaPins_Fpga_CPU_inc_pc_a1,
             FpgaPins_Fpga_CPU_inc_pc_a2,
             FpgaPins_Fpga_CPU_inc_pc_a3;

// For /fpga_pins/fpga|cpu$instr.
logic [31:0] FpgaPins_Fpga_CPU_instr_a0,
             FpgaPins_Fpga_CPU_instr_a1;

// For /fpga_pins/fpga|cpu$is_add.
logic FpgaPins_Fpga_CPU_is_add_a1;

// For /fpga_pins/fpga|cpu$is_add_op.
logic FpgaPins_Fpga_CPU_is_add_op_a1,
      FpgaPins_Fpga_CPU_is_add_op_a2,
      FpgaPins_Fpga_CPU_is_add_op_a3;

// For /fpga_pins/fpga|cpu$is_addi.
logic FpgaPins_Fpga_CPU_is_addi_a1;

// For /fpga_pins/fpga|cpu$is_and.
logic FpgaPins_Fpga_CPU_is_and_a1;

// For /fpga_pins/fpga|cpu$is_and_op.
logic FpgaPins_Fpga_CPU_is_and_op_a1,
      FpgaPins_Fpga_CPU_is_and_op_a2,
      FpgaPins_Fpga_CPU_is_and_op_a3;

// For /fpga_pins/fpga|cpu$is_andi.
logic FpgaPins_Fpga_CPU_is_andi_a1;

// For /fpga_pins/fpga|cpu$is_auipc.
logic FpgaPins_Fpga_CPU_is_auipc_a1,
      FpgaPins_Fpga_CPU_is_auipc_a2;

// For /fpga_pins/fpga|cpu$is_b_instr.
logic FpgaPins_Fpga_CPU_is_b_instr_a1,
      FpgaPins_Fpga_CPU_is_b_instr_a2;

// For /fpga_pins/fpga|cpu$is_beq.
logic FpgaPins_Fpga_CPU_is_beq_a1,
      FpgaPins_Fpga_CPU_is_beq_a2,
      FpgaPins_Fpga_CPU_is_beq_a3;

// For /fpga_pins/fpga|cpu$is_bge.
logic FpgaPins_Fpga_CPU_is_bge_a1,
      FpgaPins_Fpga_CPU_is_bge_a2,
      FpgaPins_Fpga_CPU_is_bge_a3;

// For /fpga_pins/fpga|cpu$is_bgeu.
logic FpgaPins_Fpga_CPU_is_bgeu_a1,
      FpgaPins_Fpga_CPU_is_bgeu_a2,
      FpgaPins_Fpga_CPU_is_bgeu_a3;

// For /fpga_pins/fpga|cpu$is_blt.
logic FpgaPins_Fpga_CPU_is_blt_a1,
      FpgaPins_Fpga_CPU_is_blt_a2,
      FpgaPins_Fpga_CPU_is_blt_a3;

// For /fpga_pins/fpga|cpu$is_bltu.
logic FpgaPins_Fpga_CPU_is_bltu_a1,
      FpgaPins_Fpga_CPU_is_bltu_a2,
      FpgaPins_Fpga_CPU_is_bltu_a3;

// For /fpga_pins/fpga|cpu$is_bne.
logic FpgaPins_Fpga_CPU_is_bne_a1,
      FpgaPins_Fpga_CPU_is_bne_a2,
      FpgaPins_Fpga_CPU_is_bne_a3;

// For /fpga_pins/fpga|cpu$is_i_instr.
logic FpgaPins_Fpga_CPU_is_i_instr_a1;

// For /fpga_pins/fpga|cpu$is_j_instr.
logic FpgaPins_Fpga_CPU_is_j_instr_a1;

// For /fpga_pins/fpga|cpu$is_jal.
logic FpgaPins_Fpga_CPU_is_jal_a1;

// For /fpga_pins/fpga|cpu$is_jalr.
logic FpgaPins_Fpga_CPU_is_jalr_a1,
      FpgaPins_Fpga_CPU_is_jalr_a2;

// For /fpga_pins/fpga|cpu$is_jump.
logic FpgaPins_Fpga_CPU_is_jump_a1,
      FpgaPins_Fpga_CPU_is_jump_a2,
      FpgaPins_Fpga_CPU_is_jump_a3;

// For /fpga_pins/fpga|cpu$is_lb.
logic FpgaPins_Fpga_CPU_is_lb_a1;

// For /fpga_pins/fpga|cpu$is_lbu.
logic FpgaPins_Fpga_CPU_is_lbu_a1;

// For /fpga_pins/fpga|cpu$is_lh.
logic FpgaPins_Fpga_CPU_is_lh_a1;

// For /fpga_pins/fpga|cpu$is_lhu.
logic FpgaPins_Fpga_CPU_is_lhu_a1;

// For /fpga_pins/fpga|cpu$is_load.
logic FpgaPins_Fpga_CPU_is_load_a1,
      FpgaPins_Fpga_CPU_is_load_a2,
      FpgaPins_Fpga_CPU_is_load_a3;

// For /fpga_pins/fpga|cpu$is_lui.
logic FpgaPins_Fpga_CPU_is_lui_a1,
      FpgaPins_Fpga_CPU_is_lui_a2,
      FpgaPins_Fpga_CPU_is_lui_a3;

// For /fpga_pins/fpga|cpu$is_lw.
logic FpgaPins_Fpga_CPU_is_lw_a1;

// For /fpga_pins/fpga|cpu$is_or.
logic FpgaPins_Fpga_CPU_is_or_a1;

// For /fpga_pins/fpga|cpu$is_or_op.
logic FpgaPins_Fpga_CPU_is_or_op_a1,
      FpgaPins_Fpga_CPU_is_or_op_a2,
      FpgaPins_Fpga_CPU_is_or_op_a3;

// For /fpga_pins/fpga|cpu$is_ori.
logic FpgaPins_Fpga_CPU_is_ori_a1;

// For /fpga_pins/fpga|cpu$is_r_instr.
logic FpgaPins_Fpga_CPU_is_r_instr_a1,
      FpgaPins_Fpga_CPU_is_r_instr_a2;

// For /fpga_pins/fpga|cpu$is_s_instr.
logic FpgaPins_Fpga_CPU_is_s_instr_a1;

// For /fpga_pins/fpga|cpu$is_sb.
logic FpgaPins_Fpga_CPU_is_sb_a1;

// For /fpga_pins/fpga|cpu$is_sh.
logic FpgaPins_Fpga_CPU_is_sh_a1;

// For /fpga_pins/fpga|cpu$is_sll.
logic FpgaPins_Fpga_CPU_is_sll_a1;

// For /fpga_pins/fpga|cpu$is_sll_op.
logic FpgaPins_Fpga_CPU_is_sll_op_a1,
      FpgaPins_Fpga_CPU_is_sll_op_a2,
      FpgaPins_Fpga_CPU_is_sll_op_a3;

// For /fpga_pins/fpga|cpu$is_slli.
logic FpgaPins_Fpga_CPU_is_slli_a1;

// For /fpga_pins/fpga|cpu$is_slt.
logic FpgaPins_Fpga_CPU_is_slt_a1;

// For /fpga_pins/fpga|cpu$is_slt_op.
logic FpgaPins_Fpga_CPU_is_slt_op_a1,
      FpgaPins_Fpga_CPU_is_slt_op_a2,
      FpgaPins_Fpga_CPU_is_slt_op_a3;

// For /fpga_pins/fpga|cpu$is_slti.
logic FpgaPins_Fpga_CPU_is_slti_a1;

// For /fpga_pins/fpga|cpu$is_sltiu.
logic FpgaPins_Fpga_CPU_is_sltiu_a1;

// For /fpga_pins/fpga|cpu$is_sltu.
logic FpgaPins_Fpga_CPU_is_sltu_a1;

// For /fpga_pins/fpga|cpu$is_sltu_op.
logic FpgaPins_Fpga_CPU_is_sltu_op_a1,
      FpgaPins_Fpga_CPU_is_sltu_op_a2,
      FpgaPins_Fpga_CPU_is_sltu_op_a3;

// For /fpga_pins/fpga|cpu$is_sra.
logic FpgaPins_Fpga_CPU_is_sra_a1;

// For /fpga_pins/fpga|cpu$is_sra_op.
logic FpgaPins_Fpga_CPU_is_sra_op_a1,
      FpgaPins_Fpga_CPU_is_sra_op_a2,
      FpgaPins_Fpga_CPU_is_sra_op_a3;

// For /fpga_pins/fpga|cpu$is_srai.
logic FpgaPins_Fpga_CPU_is_srai_a1;

// For /fpga_pins/fpga|cpu$is_srl.
logic FpgaPins_Fpga_CPU_is_srl_a1;

// For /fpga_pins/fpga|cpu$is_srl_op.
logic FpgaPins_Fpga_CPU_is_srl_op_a1,
      FpgaPins_Fpga_CPU_is_srl_op_a2,
      FpgaPins_Fpga_CPU_is_srl_op_a3;

// For /fpga_pins/fpga|cpu$is_srli.
logic FpgaPins_Fpga_CPU_is_srli_a1;

// For /fpga_pins/fpga|cpu$is_store.
logic FpgaPins_Fpga_CPU_is_store_a1,
      FpgaPins_Fpga_CPU_is_store_a2,
      FpgaPins_Fpga_CPU_is_store_a3;

// For /fpga_pins/fpga|cpu$is_sub.
logic FpgaPins_Fpga_CPU_is_sub_a1,
      FpgaPins_Fpga_CPU_is_sub_a2,
      FpgaPins_Fpga_CPU_is_sub_a3;

// For /fpga_pins/fpga|cpu$is_sw.
logic FpgaPins_Fpga_CPU_is_sw_a1;

// For /fpga_pins/fpga|cpu$is_u_instr.
logic FpgaPins_Fpga_CPU_is_u_instr_a1;

// For /fpga_pins/fpga|cpu$is_xor.
logic FpgaPins_Fpga_CPU_is_xor_a1;

// For /fpga_pins/fpga|cpu$is_xor_op.
logic FpgaPins_Fpga_CPU_is_xor_op_a1,
      FpgaPins_Fpga_CPU_is_xor_op_a2,
      FpgaPins_Fpga_CPU_is_xor_op_a3;

// For /fpga_pins/fpga|cpu$is_xori.
logic FpgaPins_Fpga_CPU_is_xori_a1;

// For /fpga_pins/fpga|cpu$ld_data.
logic [31:0] FpgaPins_Fpga_CPU_ld_data_a4,
             FpgaPins_Fpga_CPU_ld_data_a5;

// For /fpga_pins/fpga|cpu$opcode.
logic [6:0] FpgaPins_Fpga_CPU_opcode_a1;

// For /fpga_pins/fpga|cpu$pc.
logic [31:0] FpgaPins_Fpga_CPU_pc_a0,
             FpgaPins_Fpga_CPU_pc_a1,
             FpgaPins_Fpga_CPU_pc_a2;

// For /fpga_pins/fpga|cpu$rd.
logic [4:0] FpgaPins_Fpga_CPU_rd_a1,
            FpgaPins_Fpga_CPU_rd_a2,
            FpgaPins_Fpga_CPU_rd_a3,
            FpgaPins_Fpga_CPU_rd_a4,
            FpgaPins_Fpga_CPU_rd_a5;

// For /fpga_pins/fpga|cpu$rd_valid.
logic FpgaPins_Fpga_CPU_rd_valid_a1,
      FpgaPins_Fpga_CPU_rd_valid_a2,
      FpgaPins_Fpga_CPU_rd_valid_a3;

// For /fpga_pins/fpga|cpu$reset.
logic FpgaPins_Fpga_CPU_reset_a0,
      FpgaPins_Fpga_CPU_reset_a1,
      FpgaPins_Fpga_CPU_reset_a2,
      FpgaPins_Fpga_CPU_reset_a3;

// For /fpga_pins/fpga|cpu$result.
logic [31:0] FpgaPins_Fpga_CPU_result_a3;
logic [31:2] FpgaPins_Fpga_CPU_result_a4;

// For /fpga_pins/fpga|cpu$rf_rd_data1.
logic [31:0] FpgaPins_Fpga_CPU_rf_rd_data1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_data2.
logic [31:0] FpgaPins_Fpga_CPU_rf_rd_data2_a2;

// For /fpga_pins/fpga|cpu$rf_rd_en1.
logic FpgaPins_Fpga_CPU_rf_rd_en1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_en2.
logic FpgaPins_Fpga_CPU_rf_rd_en2_a2;

// For /fpga_pins/fpga|cpu$rf_rd_index1.
logic [4:0] FpgaPins_Fpga_CPU_rf_rd_index1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_index2.
logic [4:0] FpgaPins_Fpga_CPU_rf_rd_index2_a2;

// For /fpga_pins/fpga|cpu$rf_wr_data.
logic [31:0] FpgaPins_Fpga_CPU_rf_wr_data_a3;

// For /fpga_pins/fpga|cpu$rf_wr_en.
logic FpgaPins_Fpga_CPU_rf_wr_en_a3;

// For /fpga_pins/fpga|cpu$rf_wr_index.
logic [4:0] FpgaPins_Fpga_CPU_rf_wr_index_a3;

// For /fpga_pins/fpga|cpu$rs1.
logic [4:0] FpgaPins_Fpga_CPU_rs1_a1,
            FpgaPins_Fpga_CPU_rs1_a2;

// For /fpga_pins/fpga|cpu$rs1_valid.
logic FpgaPins_Fpga_CPU_rs1_valid_a1,
      FpgaPins_Fpga_CPU_rs1_valid_a2;

// For /fpga_pins/fpga|cpu$rs2.
logic [4:0] FpgaPins_Fpga_CPU_rs2_a1,
            FpgaPins_Fpga_CPU_rs2_a2;

// For /fpga_pins/fpga|cpu$rs2_valid.
logic FpgaPins_Fpga_CPU_rs2_valid_a1,
      FpgaPins_Fpga_CPU_rs2_valid_a2;

// For /fpga_pins/fpga|cpu$sltu_result.
logic [31:0] FpgaPins_Fpga_CPU_sltu_result_a3;

// For /fpga_pins/fpga|cpu$sra_result.
logic [63:0] FpgaPins_Fpga_CPU_sra_result_a3;

// For /fpga_pins/fpga|cpu$src1_value.
logic [31:0] FpgaPins_Fpga_CPU_src1_value_a2;

// For /fpga_pins/fpga|cpu$src2_value.
logic [31:0] FpgaPins_Fpga_CPU_src2_value_a2,
             FpgaPins_Fpga_CPU_src2_value_a3,
             FpgaPins_Fpga_CPU_src2_value_a4;

// For /fpga_pins/fpga|cpu$tgt_pc.
logic [31:0] FpgaPins_Fpga_CPU_tgt_pc_a3;

// For /fpga_pins/fpga|cpu$tgt_pc_op1.
logic [31:0] FpgaPins_Fpga_CPU_tgt_pc_op1_a2,
             FpgaPins_Fpga_CPU_tgt_pc_op1_a3;

// For /fpga_pins/fpga|cpu$tgt_pc_op2.
logic [31:0] FpgaPins_Fpga_CPU_tgt_pc_op2_a2,
             FpgaPins_Fpga_CPU_tgt_pc_op2_a3;

// For /fpga_pins/fpga|cpu$valid.
logic FpgaPins_Fpga_CPU_valid_a3;

// For /fpga_pins/fpga|cpu$valid_jump.
logic FpgaPins_Fpga_CPU_valid_jump_a3,
      FpgaPins_Fpga_CPU_valid_jump_a4,
      FpgaPins_Fpga_CPU_valid_jump_a5;

// For /fpga_pins/fpga|cpu$valid_load.
logic FpgaPins_Fpga_CPU_valid_load_a3,
      FpgaPins_Fpga_CPU_valid_load_a4,
      FpgaPins_Fpga_CPU_valid_load_a5;

// For /fpga_pins/fpga|cpu$valid_store.
logic FpgaPins_Fpga_CPU_valid_store_a3,
      FpgaPins_Fpga_CPU_valid_store_a4;

// For /fpga_pins/fpga|cpu$valid_taken_br.
logic FpgaPins_Fpga_CPU_valid_taken_br_a3,
      FpgaPins_Fpga_CPU_valid_taken_br_a4,
      FpgaPins_Fpga_CPU_valid_taken_br_a5;

// For /fpga_pins/fpga|cpu$valid_tgt_pc.
logic FpgaPins_Fpga_CPU_valid_tgt_pc_a3;

// For /fpga_pins/fpga|cpu/xreg$value.
logic [31:0] FpgaPins_Fpga_CPU_Xreg_value_a3 [15:0],
             FpgaPins_Fpga_CPU_Xreg_value_a4 [15:0];




   //
   // Scope: /fpga_pins
   //


      //
      // Scope: /fpga
      //


         //
         // Scope: |cpu
         //

            // Staging of $alu_op1.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_alu_op1_a3[31:0] <= FpgaPins_Fpga_CPU_alu_op1_a2[31:0];

            // Staging of $alu_op2.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_alu_op2_a3[31:0] <= FpgaPins_Fpga_CPU_alu_op2_a2[31:0];

            // Staging of $imm.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_imm_a2[31:0] <= FpgaPins_Fpga_CPU_imm_a1[31:0];

            // Staging of $inc_pc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_inc_pc_a2[31:0] <= FpgaPins_Fpga_CPU_inc_pc_a1[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_inc_pc_a3[31:0] <= FpgaPins_Fpga_CPU_inc_pc_a2[31:0];

            // Staging of $instr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_instr_a1[31:0] <= FpgaPins_Fpga_CPU_instr_a0[31:0];

            // Staging of $is_add_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_add_op_a2 <= FpgaPins_Fpga_CPU_is_add_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_add_op_a3 <= FpgaPins_Fpga_CPU_is_add_op_a2;

            // Staging of $is_and_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_and_op_a2 <= FpgaPins_Fpga_CPU_is_and_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_and_op_a3 <= FpgaPins_Fpga_CPU_is_and_op_a2;

            // Staging of $is_auipc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_auipc_a2 <= FpgaPins_Fpga_CPU_is_auipc_a1;

            // Staging of $is_b_instr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_b_instr_a2 <= FpgaPins_Fpga_CPU_is_b_instr_a1;

            // Staging of $is_beq.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_beq_a2 <= FpgaPins_Fpga_CPU_is_beq_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_beq_a3 <= FpgaPins_Fpga_CPU_is_beq_a2;

            // Staging of $is_bge.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bge_a2 <= FpgaPins_Fpga_CPU_is_bge_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bge_a3 <= FpgaPins_Fpga_CPU_is_bge_a2;

            // Staging of $is_bgeu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bgeu_a2 <= FpgaPins_Fpga_CPU_is_bgeu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bgeu_a3 <= FpgaPins_Fpga_CPU_is_bgeu_a2;

            // Staging of $is_blt.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_blt_a2 <= FpgaPins_Fpga_CPU_is_blt_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_blt_a3 <= FpgaPins_Fpga_CPU_is_blt_a2;

            // Staging of $is_bltu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bltu_a2 <= FpgaPins_Fpga_CPU_is_bltu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bltu_a3 <= FpgaPins_Fpga_CPU_is_bltu_a2;

            // Staging of $is_bne.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bne_a2 <= FpgaPins_Fpga_CPU_is_bne_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bne_a3 <= FpgaPins_Fpga_CPU_is_bne_a2;

            // Staging of $is_jalr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jalr_a2 <= FpgaPins_Fpga_CPU_is_jalr_a1;

            // Staging of $is_jump.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jump_a2 <= FpgaPins_Fpga_CPU_is_jump_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jump_a3 <= FpgaPins_Fpga_CPU_is_jump_a2;

            // Staging of $is_load.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_load_a2 <= FpgaPins_Fpga_CPU_is_load_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_load_a3 <= FpgaPins_Fpga_CPU_is_load_a2;

            // Staging of $is_lui.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_lui_a2 <= FpgaPins_Fpga_CPU_is_lui_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_lui_a3 <= FpgaPins_Fpga_CPU_is_lui_a2;

            // Staging of $is_or_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_or_op_a2 <= FpgaPins_Fpga_CPU_is_or_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_or_op_a3 <= FpgaPins_Fpga_CPU_is_or_op_a2;

            // Staging of $is_r_instr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_r_instr_a2 <= FpgaPins_Fpga_CPU_is_r_instr_a1;

            // Staging of $is_sll_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sll_op_a2 <= FpgaPins_Fpga_CPU_is_sll_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sll_op_a3 <= FpgaPins_Fpga_CPU_is_sll_op_a2;

            // Staging of $is_slt_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slt_op_a2 <= FpgaPins_Fpga_CPU_is_slt_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slt_op_a3 <= FpgaPins_Fpga_CPU_is_slt_op_a2;

            // Staging of $is_sltu_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltu_op_a2 <= FpgaPins_Fpga_CPU_is_sltu_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltu_op_a3 <= FpgaPins_Fpga_CPU_is_sltu_op_a2;

            // Staging of $is_sra_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sra_op_a2 <= FpgaPins_Fpga_CPU_is_sra_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sra_op_a3 <= FpgaPins_Fpga_CPU_is_sra_op_a2;

            // Staging of $is_srl_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srl_op_a2 <= FpgaPins_Fpga_CPU_is_srl_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srl_op_a3 <= FpgaPins_Fpga_CPU_is_srl_op_a2;

            // Staging of $is_store.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_store_a2 <= FpgaPins_Fpga_CPU_is_store_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_store_a3 <= FpgaPins_Fpga_CPU_is_store_a2;

            // Staging of $is_sub.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sub_a2 <= FpgaPins_Fpga_CPU_is_sub_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sub_a3 <= FpgaPins_Fpga_CPU_is_sub_a2;

            // Staging of $is_xor_op.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xor_op_a2 <= FpgaPins_Fpga_CPU_is_xor_op_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xor_op_a3 <= FpgaPins_Fpga_CPU_is_xor_op_a2;

            // Staging of $ld_data.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_ld_data_a5[31:0] <= FpgaPins_Fpga_CPU_ld_data_a4[31:0];

            // Staging of $pc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_pc_a1[31:0] <= FpgaPins_Fpga_CPU_pc_a0[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_pc_a2[31:0] <= FpgaPins_Fpga_CPU_pc_a1[31:0];

            // Staging of $rd.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a2[4:0] <= FpgaPins_Fpga_CPU_rd_a1[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a3[4:0] <= FpgaPins_Fpga_CPU_rd_a2[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a4[4:0] <= FpgaPins_Fpga_CPU_rd_a3[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a5[4:0] <= FpgaPins_Fpga_CPU_rd_a4[4:0];

            // Staging of $rd_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_valid_a2 <= FpgaPins_Fpga_CPU_rd_valid_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_valid_a3 <= FpgaPins_Fpga_CPU_rd_valid_a2;

            // Staging of $reset.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a1 <= FpgaPins_Fpga_CPU_reset_a0;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a2 <= FpgaPins_Fpga_CPU_reset_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a3 <= FpgaPins_Fpga_CPU_reset_a2;

            // Staging of $result.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_result_a4[31:2] <= FpgaPins_Fpga_CPU_result_a3[31:2];

            // Staging of $rs1.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs1_a2[4:0] <= FpgaPins_Fpga_CPU_rs1_a1[4:0];

            // Staging of $rs1_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs1_valid_a2 <= FpgaPins_Fpga_CPU_rs1_valid_a1;

            // Staging of $rs2.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs2_a2[4:0] <= FpgaPins_Fpga_CPU_rs2_a1[4:0];

            // Staging of $rs2_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs2_valid_a2 <= FpgaPins_Fpga_CPU_rs2_valid_a1;

            // Staging of $src2_value.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_src2_value_a3[31:0] <= FpgaPins_Fpga_CPU_src2_value_a2[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_src2_value_a4[31:0] <= FpgaPins_Fpga_CPU_src2_value_a3[31:0];

            // Staging of $tgt_pc_op1.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_tgt_pc_op1_a3[31:0] <= FpgaPins_Fpga_CPU_tgt_pc_op1_a2[31:0];

            // Staging of $tgt_pc_op2.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_tgt_pc_op2_a3[31:0] <= FpgaPins_Fpga_CPU_tgt_pc_op2_a2[31:0];

            // Staging of $valid_jump.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_jump_a4 <= FpgaPins_Fpga_CPU_valid_jump_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_jump_a5 <= FpgaPins_Fpga_CPU_valid_jump_a4;

            // Staging of $valid_load.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_load_a4 <= FpgaPins_Fpga_CPU_valid_load_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_load_a5 <= FpgaPins_Fpga_CPU_valid_load_a4;

            // Staging of $valid_store.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_store_a4 <= FpgaPins_Fpga_CPU_valid_store_a3;

            // Staging of $valid_taken_br.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_taken_br_a4 <= FpgaPins_Fpga_CPU_valid_taken_br_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_taken_br_a5 <= FpgaPins_Fpga_CPU_valid_taken_br_a4;


            //
            // Scope: /xreg[15:0]
            //
            for (xreg = 0; xreg <= 15; xreg++) begin : L1gen_FpgaPins_Fpga_CPU_Xreg
               // Staging of $value.
               always_ff @(posedge clk) FpgaPins_Fpga_CPU_Xreg_value_a4[xreg][31:0] <= FpgaPins_Fpga_CPU_Xreg_value_a3[xreg][31:0];

            end







//
// Debug Signals
//

   if (1) begin : DEBUG_SIGS_GTKWAVE

      (* keep *) logic [7:0] \@0$slideswitch ;
      assign \@0$slideswitch = L0_slideswitch_a0;
      (* keep *) logic  \@0$sseg_decimal_point_n ;
      assign \@0$sseg_decimal_point_n = L0_sseg_decimal_point_n_a0;
      (* keep *) logic [7:0] \@0$sseg_digit_n ;
      assign \@0$sseg_digit_n = L0_sseg_digit_n_a0;
      (* keep *) logic [6:0] \@0$sseg_segment_n ;
      assign \@0$sseg_segment_n = L0_sseg_segment_n_a0;

      //
      // Scope: /digit[0:0]
      //
      for (digit = 0; digit <= 0; digit++) begin : \/digit 

         //
         // Scope: /leds[7:0]
         //
         for (leds = 0; leds <= 7; leds++) begin : \/leds 
            (* keep *) logic  \//@0$viz_lit ;
            assign \//@0$viz_lit = L1_Digit[digit].L2_Leds[leds].L2_viz_lit_a0;
         end
      end

      //
      // Scope: /fpga_pins
      //
      if (1) begin : \/fpga_pins 

         //
         // Scope: /fpga
         //
         if (1) begin : \/fpga 

            //
            // Scope: |cpu
            //
            if (1) begin : P_cpu
               (* keep *) logic [31:0] \///@2$alu_op1 ;
               assign \///@2$alu_op1 = FpgaPins_Fpga_CPU_alu_op1_a2;
               (* keep *) logic [31:0] \///@2$alu_op2 ;
               assign \///@2$alu_op2 = FpgaPins_Fpga_CPU_alu_op2_a2;
               (* keep *) logic [2:0] \///@1$funct3 ;
               assign \///@1$funct3 = FpgaPins_Fpga_CPU_funct3_a1;
               (* keep *) logic [6:0] \///@1$funct7 ;
               assign \///@1$funct7 = FpgaPins_Fpga_CPU_funct7_a1;
               (* keep *) logic [31:0] \///@1$imm ;
               assign \///@1$imm = FpgaPins_Fpga_CPU_imm_a1;
               (* keep *) logic [31:0] \///@1$inc_pc ;
               assign \///@1$inc_pc = FpgaPins_Fpga_CPU_inc_pc_a1;
               (* keep *) logic [31:0] \///@0$instr ;
               assign \///@0$instr = FpgaPins_Fpga_CPU_instr_a0;
               (* keep *) logic  \///@1$is_add ;
               assign \///@1$is_add = FpgaPins_Fpga_CPU_is_add_a1;
               (* keep *) logic  \///@1$is_add_op ;
               assign \///@1$is_add_op = FpgaPins_Fpga_CPU_is_add_op_a1;
               (* keep *) logic  \///@1$is_addi ;
               assign \///@1$is_addi = FpgaPins_Fpga_CPU_is_addi_a1;
               (* keep *) logic  \///@1$is_and ;
               assign \///@1$is_and = FpgaPins_Fpga_CPU_is_and_a1;
               (* keep *) logic  \///@1$is_and_op ;
               assign \///@1$is_and_op = FpgaPins_Fpga_CPU_is_and_op_a1;
               (* keep *) logic  \///@1$is_andi ;
               assign \///@1$is_andi = FpgaPins_Fpga_CPU_is_andi_a1;
               (* keep *) logic  \///@1$is_auipc ;
               assign \///@1$is_auipc = FpgaPins_Fpga_CPU_is_auipc_a1;
               (* keep *) logic  \///@1$is_b_instr ;
               assign \///@1$is_b_instr = FpgaPins_Fpga_CPU_is_b_instr_a1;
               (* keep *) logic  \///@1$is_beq ;
               assign \///@1$is_beq = FpgaPins_Fpga_CPU_is_beq_a1;
               (* keep *) logic  \///@1$is_bge ;
               assign \///@1$is_bge = FpgaPins_Fpga_CPU_is_bge_a1;
               (* keep *) logic  \///@1$is_bgeu ;
               assign \///@1$is_bgeu = FpgaPins_Fpga_CPU_is_bgeu_a1;
               (* keep *) logic  \///@1$is_blt ;
               assign \///@1$is_blt = FpgaPins_Fpga_CPU_is_blt_a1;
               (* keep *) logic  \///@1$is_bltu ;
               assign \///@1$is_bltu = FpgaPins_Fpga_CPU_is_bltu_a1;
               (* keep *) logic  \///@1$is_bne ;
               assign \///@1$is_bne = FpgaPins_Fpga_CPU_is_bne_a1;
               (* keep *) logic  \///@1$is_i_instr ;
               assign \///@1$is_i_instr = FpgaPins_Fpga_CPU_is_i_instr_a1;
               (* keep *) logic  \///@1$is_j_instr ;
               assign \///@1$is_j_instr = FpgaPins_Fpga_CPU_is_j_instr_a1;
               (* keep *) logic  \///@1$is_jal ;
               assign \///@1$is_jal = FpgaPins_Fpga_CPU_is_jal_a1;
               (* keep *) logic  \///@1$is_jalr ;
               assign \///@1$is_jalr = FpgaPins_Fpga_CPU_is_jalr_a1;
               (* keep *) logic  \///@1$is_jump ;
               assign \///@1$is_jump = FpgaPins_Fpga_CPU_is_jump_a1;
               (* keep *) logic  \///@1$is_lb ;
               assign \///@1$is_lb = FpgaPins_Fpga_CPU_is_lb_a1;
               (* keep *) logic  \///@1$is_lbu ;
               assign \///@1$is_lbu = FpgaPins_Fpga_CPU_is_lbu_a1;
               (* keep *) logic  \///@1$is_lh ;
               assign \///@1$is_lh = FpgaPins_Fpga_CPU_is_lh_a1;
               (* keep *) logic  \///@1$is_lhu ;
               assign \///@1$is_lhu = FpgaPins_Fpga_CPU_is_lhu_a1;
               (* keep *) logic  \///@1$is_load ;
               assign \///@1$is_load = FpgaPins_Fpga_CPU_is_load_a1;
               (* keep *) logic  \///@1$is_lui ;
               assign \///@1$is_lui = FpgaPins_Fpga_CPU_is_lui_a1;
               (* keep *) logic  \///@1$is_lw ;
               assign \///@1$is_lw = FpgaPins_Fpga_CPU_is_lw_a1;
               (* keep *) logic  \///@1$is_or ;
               assign \///@1$is_or = FpgaPins_Fpga_CPU_is_or_a1;
               (* keep *) logic  \///@1$is_or_op ;
               assign \///@1$is_or_op = FpgaPins_Fpga_CPU_is_or_op_a1;
               (* keep *) logic  \///@1$is_ori ;
               assign \///@1$is_ori = FpgaPins_Fpga_CPU_is_ori_a1;
               (* keep *) logic  \///@1$is_r_instr ;
               assign \///@1$is_r_instr = FpgaPins_Fpga_CPU_is_r_instr_a1;
               (* keep *) logic  \///@1$is_s_instr ;
               assign \///@1$is_s_instr = FpgaPins_Fpga_CPU_is_s_instr_a1;
               (* keep *) logic  \///@1$is_sb ;
               assign \///@1$is_sb = FpgaPins_Fpga_CPU_is_sb_a1;
               (* keep *) logic  \///@1$is_sh ;
               assign \///@1$is_sh = FpgaPins_Fpga_CPU_is_sh_a1;
               (* keep *) logic  \///@1$is_sll ;
               assign \///@1$is_sll = FpgaPins_Fpga_CPU_is_sll_a1;
               (* keep *) logic  \///@1$is_sll_op ;
               assign \///@1$is_sll_op = FpgaPins_Fpga_CPU_is_sll_op_a1;
               (* keep *) logic  \///@1$is_slli ;
               assign \///@1$is_slli = FpgaPins_Fpga_CPU_is_slli_a1;
               (* keep *) logic  \///@1$is_slt ;
               assign \///@1$is_slt = FpgaPins_Fpga_CPU_is_slt_a1;
               (* keep *) logic  \///@1$is_slt_op ;
               assign \///@1$is_slt_op = FpgaPins_Fpga_CPU_is_slt_op_a1;
               (* keep *) logic  \///@1$is_slti ;
               assign \///@1$is_slti = FpgaPins_Fpga_CPU_is_slti_a1;
               (* keep *) logic  \///@1$is_sltiu ;
               assign \///@1$is_sltiu = FpgaPins_Fpga_CPU_is_sltiu_a1;
               (* keep *) logic  \///@1$is_sltu ;
               assign \///@1$is_sltu = FpgaPins_Fpga_CPU_is_sltu_a1;
               (* keep *) logic  \///@1$is_sltu_op ;
               assign \///@1$is_sltu_op = FpgaPins_Fpga_CPU_is_sltu_op_a1;
               (* keep *) logic  \///@1$is_sra ;
               assign \///@1$is_sra = FpgaPins_Fpga_CPU_is_sra_a1;
               (* keep *) logic  \///@1$is_sra_op ;
               assign \///@1$is_sra_op = FpgaPins_Fpga_CPU_is_sra_op_a1;
               (* keep *) logic  \///@1$is_srai ;
               assign \///@1$is_srai = FpgaPins_Fpga_CPU_is_srai_a1;
               (* keep *) logic  \///@1$is_srl ;
               assign \///@1$is_srl = FpgaPins_Fpga_CPU_is_srl_a1;
               (* keep *) logic  \///@1$is_srl_op ;
               assign \///@1$is_srl_op = FpgaPins_Fpga_CPU_is_srl_op_a1;
               (* keep *) logic  \///@1$is_srli ;
               assign \///@1$is_srli = FpgaPins_Fpga_CPU_is_srli_a1;
               (* keep *) logic  \///@1$is_store ;
               assign \///@1$is_store = FpgaPins_Fpga_CPU_is_store_a1;
               (* keep *) logic  \///@1$is_sub ;
               assign \///@1$is_sub = FpgaPins_Fpga_CPU_is_sub_a1;
               (* keep *) logic  \///@1$is_sw ;
               assign \///@1$is_sw = FpgaPins_Fpga_CPU_is_sw_a1;
               (* keep *) logic  \///@1$is_u_instr ;
               assign \///@1$is_u_instr = FpgaPins_Fpga_CPU_is_u_instr_a1;
               (* keep *) logic  \///@1$is_xor ;
               assign \///@1$is_xor = FpgaPins_Fpga_CPU_is_xor_a1;
               (* keep *) logic  \///@1$is_xor_op ;
               assign \///@1$is_xor_op = FpgaPins_Fpga_CPU_is_xor_op_a1;
               (* keep *) logic  \///@1$is_xori ;
               assign \///@1$is_xori = FpgaPins_Fpga_CPU_is_xori_a1;
               (* keep *) logic [31:0] \///@4$ld_data ;
               assign \///@4$ld_data = FpgaPins_Fpga_CPU_ld_data_a4;
               (* keep *) logic [6:0] \///@1$opcode ;
               assign \///@1$opcode = FpgaPins_Fpga_CPU_opcode_a1;
               (* keep *) logic [31:0] \///@0$pc ;
               assign \///@0$pc = FpgaPins_Fpga_CPU_pc_a0;
               (* keep *) logic [4:0] \///@1$rd ;
               assign \///@1$rd = FpgaPins_Fpga_CPU_rd_a1;
               (* keep *) logic  \///@1$rd_valid ;
               assign \///@1$rd_valid = FpgaPins_Fpga_CPU_rd_valid_a1;
               (* keep *) logic  \///@0$reset ;
               assign \///@0$reset = FpgaPins_Fpga_CPU_reset_a0;
               (* keep *) logic [31:0] \///@3$result ;
               assign \///@3$result = FpgaPins_Fpga_CPU_result_a3;
               (* keep *) logic [31:0] \///?$rf_rd_en1@2$rf_rd_data1 ;
               assign \///?$rf_rd_en1@2$rf_rd_data1 = FpgaPins_Fpga_CPU_rf_rd_data1_a2;
               (* keep *) logic [31:0] \///?$rf_rd_en2@2$rf_rd_data2 ;
               assign \///?$rf_rd_en2@2$rf_rd_data2 = FpgaPins_Fpga_CPU_rf_rd_data2_a2;
               (* keep *) logic  \///@2$rf_rd_en1 ;
               assign \///@2$rf_rd_en1 = FpgaPins_Fpga_CPU_rf_rd_en1_a2;
               (* keep *) logic  \///@2$rf_rd_en2 ;
               assign \///@2$rf_rd_en2 = FpgaPins_Fpga_CPU_rf_rd_en2_a2;
               (* keep *) logic [4:0] \///@2$rf_rd_index1 ;
               assign \///@2$rf_rd_index1 = FpgaPins_Fpga_CPU_rf_rd_index1_a2;
               (* keep *) logic [4:0] \///@2$rf_rd_index2 ;
               assign \///@2$rf_rd_index2 = FpgaPins_Fpga_CPU_rf_rd_index2_a2;
               (* keep *) logic [31:0] \///@3$rf_wr_data ;
               assign \///@3$rf_wr_data = FpgaPins_Fpga_CPU_rf_wr_data_a3;
               (* keep *) logic  \///@3$rf_wr_en ;
               assign \///@3$rf_wr_en = FpgaPins_Fpga_CPU_rf_wr_en_a3;
               (* keep *) logic [4:0] \///@3$rf_wr_index ;
               assign \///@3$rf_wr_index = FpgaPins_Fpga_CPU_rf_wr_index_a3;
               (* keep *) logic [4:0] \///@1$rs1 ;
               assign \///@1$rs1 = FpgaPins_Fpga_CPU_rs1_a1;
               (* keep *) logic  \///@1$rs1_valid ;
               assign \///@1$rs1_valid = FpgaPins_Fpga_CPU_rs1_valid_a1;
               (* keep *) logic [4:0] \///@1$rs2 ;
               assign \///@1$rs2 = FpgaPins_Fpga_CPU_rs2_a1;
               (* keep *) logic  \///@1$rs2_valid ;
               assign \///@1$rs2_valid = FpgaPins_Fpga_CPU_rs2_valid_a1;
               (* keep *) logic [31:0] \///@3$sltu_result ;
               assign \///@3$sltu_result = FpgaPins_Fpga_CPU_sltu_result_a3;
               (* keep *) logic [63:0] \///@3$sra_result ;
               assign \///@3$sra_result = FpgaPins_Fpga_CPU_sra_result_a3;
               (* keep *) logic [31:0] \///@2$src1_value ;
               assign \///@2$src1_value = FpgaPins_Fpga_CPU_src1_value_a2;
               (* keep *) logic [31:0] \///@2$src2_value ;
               assign \///@2$src2_value = FpgaPins_Fpga_CPU_src2_value_a2;
               (* keep *) logic [31:0] \///@3$tgt_pc ;
               assign \///@3$tgt_pc = FpgaPins_Fpga_CPU_tgt_pc_a3;
               (* keep *) logic [31:0] \///@2$tgt_pc_op1 ;
               assign \///@2$tgt_pc_op1 = FpgaPins_Fpga_CPU_tgt_pc_op1_a2;
               (* keep *) logic [31:0] \///@2$tgt_pc_op2 ;
               assign \///@2$tgt_pc_op2 = FpgaPins_Fpga_CPU_tgt_pc_op2_a2;
               (* keep *) logic  \///@3$valid ;
               assign \///@3$valid = FpgaPins_Fpga_CPU_valid_a3;
               (* keep *) logic  \///@3$valid_jump ;
               assign \///@3$valid_jump = FpgaPins_Fpga_CPU_valid_jump_a3;
               (* keep *) logic  \///@3$valid_load ;
               assign \///@3$valid_load = FpgaPins_Fpga_CPU_valid_load_a3;
               (* keep *) logic  \///@3$valid_store ;
               assign \///@3$valid_store = FpgaPins_Fpga_CPU_valid_store_a3;
               (* keep *) logic  \///@3$valid_taken_br ;
               assign \///@3$valid_taken_br = FpgaPins_Fpga_CPU_valid_taken_br_a3;
               (* keep *) logic  \///@3$valid_tgt_pc ;
               assign \///@3$valid_tgt_pc = FpgaPins_Fpga_CPU_valid_tgt_pc_a3;

               //
               // Scope: /xreg[15:0]
               //
               for (xreg = 0; xreg <= 15; xreg++) begin : \/xreg 
                  (* keep *) logic [31:0] \////@3$value ;
                  assign \////@3$value = FpgaPins_Fpga_CPU_Xreg_value_a3[xreg];
                  (* keep *) logic  \////@3$wr ;
                  assign \////@3$wr = L1_FpgaPins_Fpga_CPU_Xreg[xreg].L1_wr_a3;
               end
            end
         end
      end

      //
      // Scope: /switch[7:0]
      //
      for (switch = 0; switch <= 7; switch++) begin : \/switch 
         (* keep *) logic  \/@0$viz_switch ;
         assign \/@0$viz_switch = L1_Switch[switch].L1_viz_switch_a0;
      end


   end

// ---------- Generated Code Ends ----------
//_\TLV
   /* verilator lint_off UNOPTFLAT */
   // Connect Tiny Tapeout I/Os to Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/35e36bd144fddd75495d4cbc01c4fc50ac5bde6f/tlvlib/tinytapeoutlib.tlv 76   // Instantiated from top.tlv, 400 as: m5+tt_connections()
      assign L0_slideswitch_a0[7:0] = ui_in;
      assign L0_sseg_segment_n_a0[6:0] = ~ uo_out[6:0];
      assign L0_sseg_decimal_point_n_a0 = ~ uo_out[7];
      assign L0_sseg_digit_n_a0[7:0] = 8'b11111110;
   //_\end_source

   // Instantiate the Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 307   // Instantiated from top.tlv, 403 as: m5+board(/top, /fpga, 7, $, , cpu)
      
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 355   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 309 as: m4+thanks(m5__l(309)m5_eval(m5_get(BOARD_THANKS_ARGS)))
         //_/thanks
            
      //_\end_source
      
   
      // Board VIZ.
   
      // Board Image.
      
      //_/fpga_pins
         
         //_/fpga
            //_\source top.tlv 96   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 340 as: m4+cpu.
            
               //_\source M5-FN-riscv_gen 0   // Instantiated from top.tlv, 98 as: m5+riscv_gen()
                  
               //_\end_source
               //_\source M5-FN-riscv_sum_prog 0   // Instantiated from top.tlv, 99 as: m5+riscv_sum_prog()
                  // Inst #0: ADD x10, x0, x0
                  // Inst #1: ADD x14, x10, x0
                  // Inst #2: ADDI x12, x10, 10
                  // Inst #3: ADD x13, x10, x0
                  // Inst #4: ADD x14, x13, x14
                  // Inst #5: ADDI x13, x13, 1
                  // Inst #6: BLT x13, x12, loop
                  // Inst #7: ADD x10, x14, x0
                  // Inst #8: SW x0, x10, 4
                  // Inst #9: LW x15, x0, 4
                  // Inst #10: JALR x1, x0, 0
                  
               //_\end_source
               
               //_|cpu
                  //_@0 // Instruction Fetch, PC Select
                     assign FpgaPins_Fpga_CPU_reset_a0 = reset;
                     assign FpgaPins_Fpga_CPU_pc_a0[31:0] =
                        FpgaPins_Fpga_CPU_reset_a0             ? 32'h0000_0000 :
                        FpgaPins_Fpga_CPU_reset_a1          ? 32'h0000_0000 :
                        FpgaPins_Fpga_CPU_valid_tgt_pc_a3   ? FpgaPins_Fpga_CPU_tgt_pc_a3 :
                        FpgaPins_Fpga_CPU_valid_load_a3     ? FpgaPins_Fpga_CPU_inc_pc_a3 :
                                             FpgaPins_Fpga_CPU_inc_pc_a1;
                     assign imem_rd_en = ! (FpgaPins_Fpga_CPU_reset_a0 || FpgaPins_Fpga_CPU_reset_a1);
                     assign imem_rd_addr = FpgaPins_Fpga_CPU_pc_a0[IMEM_BYTE_ADDR_WIDTH-1:2];
                     assign FpgaPins_Fpga_CPU_instr_a0[31:0] = imem_rd_data[31:0];
            
                  //_@1 // Instruction Decode, PC Increment
                     assign FpgaPins_Fpga_CPU_inc_pc_a1[31:0] = FpgaPins_Fpga_CPU_pc_a1 + 32'h4;
            
                     // Instruction Fields
                     assign FpgaPins_Fpga_CPU_opcode_a1[6:0] = FpgaPins_Fpga_CPU_instr_a1[6:0];
                     assign FpgaPins_Fpga_CPU_funct3_a1[2:0] = FpgaPins_Fpga_CPU_instr_a1[14:12];
                     assign FpgaPins_Fpga_CPU_funct7_a1[6:0] = FpgaPins_Fpga_CPU_instr_a1[31:25];
                     assign FpgaPins_Fpga_CPU_rd_a1[4:0] = FpgaPins_Fpga_CPU_instr_a1[11:7];
                     assign FpgaPins_Fpga_CPU_rs1_a1[4:0] = FpgaPins_Fpga_CPU_instr_a1[19:15];
                     assign FpgaPins_Fpga_CPU_rs2_a1[4:0] = FpgaPins_Fpga_CPU_instr_a1[24:20];
                     assign FpgaPins_Fpga_CPU_imm_a1[31:0] =
                        FpgaPins_Fpga_CPU_is_s_instr_a1 ? {{21{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[30:25], FpgaPins_Fpga_CPU_instr_a1[11:7]} :
                        FpgaPins_Fpga_CPU_is_b_instr_a1 ? {{20{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[7], FpgaPins_Fpga_CPU_instr_a1[30:25], FpgaPins_Fpga_CPU_instr_a1[11:8], 1'b0} :
                        FpgaPins_Fpga_CPU_is_u_instr_a1 ? {FpgaPins_Fpga_CPU_instr_a1[31:12], {12{1'b0}}} :
                        FpgaPins_Fpga_CPU_is_j_instr_a1 ? {{12{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[19:12], FpgaPins_Fpga_CPU_instr_a1[20], FpgaPins_Fpga_CPU_instr_a1[30:25], FpgaPins_Fpga_CPU_instr_a1[24:21], 1'b0} :
                        //default to I-type format for simplicity
                                      {{21{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[30:20]};
            
                     // Instruction Set
                     assign FpgaPins_Fpga_CPU_is_lui_a1   = FpgaPins_Fpga_CPU_opcode_a1 == 7'b0110111;
                     assign FpgaPins_Fpga_CPU_is_auipc_a1 = FpgaPins_Fpga_CPU_opcode_a1 == 7'b0010111;
                     assign FpgaPins_Fpga_CPU_is_jal_a1   = FpgaPins_Fpga_CPU_opcode_a1 == 7'b1101111;
                     assign FpgaPins_Fpga_CPU_is_jalr_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b000_1100111;
                     assign FpgaPins_Fpga_CPU_is_beq_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b000_1100011;
                     assign FpgaPins_Fpga_CPU_is_bne_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b001_1100011;
                     assign FpgaPins_Fpga_CPU_is_blt_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b100_1100011;
                     assign FpgaPins_Fpga_CPU_is_bge_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b101_1100011;
                     assign FpgaPins_Fpga_CPU_is_bltu_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b110_1100011;
                     assign FpgaPins_Fpga_CPU_is_bgeu_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b111_1100011;
                     assign FpgaPins_Fpga_CPU_is_lb_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b000_0000011;
                     assign FpgaPins_Fpga_CPU_is_lh_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b001_0000011;
                     assign FpgaPins_Fpga_CPU_is_lw_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b010_0000011;
                     assign FpgaPins_Fpga_CPU_is_lbu_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b100_0000011;
                     assign FpgaPins_Fpga_CPU_is_lhu_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b101_0000011;
                     assign FpgaPins_Fpga_CPU_is_sb_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b000_0100011;
                     assign FpgaPins_Fpga_CPU_is_sh_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b001_0100011;
                     assign FpgaPins_Fpga_CPU_is_sw_a1    = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b010_0100011;
                     assign FpgaPins_Fpga_CPU_is_addi_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b000_0010011;
                     assign FpgaPins_Fpga_CPU_is_slti_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b010_0010011;
                     assign FpgaPins_Fpga_CPU_is_sltiu_a1 = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b011_0010011;
                     assign FpgaPins_Fpga_CPU_is_xori_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b100_0010011;
                     assign FpgaPins_Fpga_CPU_is_ori_a1   = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b110_0010011;
                     assign FpgaPins_Fpga_CPU_is_andi_a1  = {FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 10'b111_0010011;
                     assign FpgaPins_Fpga_CPU_is_slli_a1  = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_001_0010011;
                     assign FpgaPins_Fpga_CPU_is_srli_a1  = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_101_0010011;
                     assign FpgaPins_Fpga_CPU_is_srai_a1  = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0100000_101_0010011;
                     assign FpgaPins_Fpga_CPU_is_add_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_000_0110011;
                     assign FpgaPins_Fpga_CPU_is_sub_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0100000_000_0110011;
                     assign FpgaPins_Fpga_CPU_is_sll_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_001_0110011;
                     assign FpgaPins_Fpga_CPU_is_slt_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_010_0110011;
                     assign FpgaPins_Fpga_CPU_is_sltu_a1  = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_011_0110011;
                     assign FpgaPins_Fpga_CPU_is_xor_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_100_0110011;
                     assign FpgaPins_Fpga_CPU_is_srl_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_101_0110011;
                     assign FpgaPins_Fpga_CPU_is_sra_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0100000_101_0110011;
                     assign FpgaPins_Fpga_CPU_is_or_a1    = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_110_0110011;
                     assign FpgaPins_Fpga_CPU_is_and_a1   = {FpgaPins_Fpga_CPU_funct7_a1, FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1} == 17'b0000000_111_0110011;
            
                     // Instruction Categories
                     assign FpgaPins_Fpga_CPU_is_load_a1    = FpgaPins_Fpga_CPU_is_lb_a1 | FpgaPins_Fpga_CPU_is_lh_a1 | FpgaPins_Fpga_CPU_is_lw_a1 | FpgaPins_Fpga_CPU_is_lbu_a1 | FpgaPins_Fpga_CPU_is_lhu_a1;
                     assign FpgaPins_Fpga_CPU_is_store_a1   = FpgaPins_Fpga_CPU_is_sb_a1 | FpgaPins_Fpga_CPU_is_sh_a1 | FpgaPins_Fpga_CPU_is_sw_a1;
                     assign FpgaPins_Fpga_CPU_is_jump_a1    = FpgaPins_Fpga_CPU_is_jal_a1  | FpgaPins_Fpga_CPU_is_jalr_a1;
                     assign FpgaPins_Fpga_CPU_is_add_op_a1  = FpgaPins_Fpga_CPU_is_add_a1  | FpgaPins_Fpga_CPU_is_addi_a1 | FpgaPins_Fpga_CPU_is_auipc_a1 | FpgaPins_Fpga_CPU_is_jump_a1 | FpgaPins_Fpga_CPU_is_load_a1 | FpgaPins_Fpga_CPU_is_store_a1;
                     assign FpgaPins_Fpga_CPU_is_and_op_a1  = FpgaPins_Fpga_CPU_is_and_a1  | FpgaPins_Fpga_CPU_is_andi_a1;
                     assign FpgaPins_Fpga_CPU_is_or_op_a1   = FpgaPins_Fpga_CPU_is_or_a1   | FpgaPins_Fpga_CPU_is_ori_a1;
                     assign FpgaPins_Fpga_CPU_is_sll_op_a1  = FpgaPins_Fpga_CPU_is_sll_a1  | FpgaPins_Fpga_CPU_is_slli_a1;
                     assign FpgaPins_Fpga_CPU_is_slt_op_a1  = FpgaPins_Fpga_CPU_is_slt_a1  | FpgaPins_Fpga_CPU_is_slti_a1  | FpgaPins_Fpga_CPU_is_blt_a1  | FpgaPins_Fpga_CPU_is_bge_a1;
                     assign FpgaPins_Fpga_CPU_is_sltu_op_a1 = FpgaPins_Fpga_CPU_is_sltu_a1 | FpgaPins_Fpga_CPU_is_sltiu_a1 | FpgaPins_Fpga_CPU_is_bltu_a1 | FpgaPins_Fpga_CPU_is_bgeu_a1;
                     assign FpgaPins_Fpga_CPU_is_sra_op_a1  = FpgaPins_Fpga_CPU_is_sra_a1  | FpgaPins_Fpga_CPU_is_srai_a1;
                     assign FpgaPins_Fpga_CPU_is_srl_op_a1  = FpgaPins_Fpga_CPU_is_srl_a1  | FpgaPins_Fpga_CPU_is_srli_a1;
                     assign FpgaPins_Fpga_CPU_is_xor_op_a1  = FpgaPins_Fpga_CPU_is_xor_a1  | FpgaPins_Fpga_CPU_is_xori_a1;
            
                     // Instruction Types
                     assign FpgaPins_Fpga_CPU_is_r_instr_a1 = FpgaPins_Fpga_CPU_is_add_a1 | FpgaPins_Fpga_CPU_is_sub_a1 | FpgaPins_Fpga_CPU_is_sll_a1 | FpgaPins_Fpga_CPU_is_slt_a1 | FpgaPins_Fpga_CPU_is_sltu_a1 | FpgaPins_Fpga_CPU_is_xor_a1 | FpgaPins_Fpga_CPU_is_srl_a1 | FpgaPins_Fpga_CPU_is_sra_a1 | FpgaPins_Fpga_CPU_is_or_a1 | FpgaPins_Fpga_CPU_is_and_a1;
                     assign FpgaPins_Fpga_CPU_is_i_instr_a1 = FpgaPins_Fpga_CPU_is_jalr_a1 | FpgaPins_Fpga_CPU_is_load_a1 | FpgaPins_Fpga_CPU_is_addi_a1 | FpgaPins_Fpga_CPU_is_slti_a1 | FpgaPins_Fpga_CPU_is_sltiu_a1 | FpgaPins_Fpga_CPU_is_xori_a1 | FpgaPins_Fpga_CPU_is_ori_a1 | FpgaPins_Fpga_CPU_is_andi_a1 | FpgaPins_Fpga_CPU_is_slli_a1 | FpgaPins_Fpga_CPU_is_srli_a1 | FpgaPins_Fpga_CPU_is_srai_a1;
                     assign FpgaPins_Fpga_CPU_is_s_instr_a1 = FpgaPins_Fpga_CPU_is_store_a1;
                     assign FpgaPins_Fpga_CPU_is_b_instr_a1 = FpgaPins_Fpga_CPU_is_beq_a1 | FpgaPins_Fpga_CPU_is_bne_a1 | FpgaPins_Fpga_CPU_is_blt_a1 | FpgaPins_Fpga_CPU_is_bge_a1 | FpgaPins_Fpga_CPU_is_bltu_a1 | FpgaPins_Fpga_CPU_is_bgeu_a1;
                     assign FpgaPins_Fpga_CPU_is_u_instr_a1 = FpgaPins_Fpga_CPU_is_lui_a1 | FpgaPins_Fpga_CPU_is_auipc_a1;
                     assign FpgaPins_Fpga_CPU_is_j_instr_a1 = FpgaPins_Fpga_CPU_is_jal_a1;
            
                     // Validity
                     assign FpgaPins_Fpga_CPU_rd_valid_a1    = !FpgaPins_Fpga_CPU_reset_a1 & (FpgaPins_Fpga_CPU_is_r_instr_a1 | FpgaPins_Fpga_CPU_is_i_instr_a1 | FpgaPins_Fpga_CPU_is_u_instr_a1 | FpgaPins_Fpga_CPU_is_j_instr_a1);
                     assign FpgaPins_Fpga_CPU_rs1_valid_a1   = !FpgaPins_Fpga_CPU_reset_a1 & (FpgaPins_Fpga_CPU_is_r_instr_a1 | FpgaPins_Fpga_CPU_is_i_instr_a1 | FpgaPins_Fpga_CPU_is_s_instr_a1 | FpgaPins_Fpga_CPU_is_b_instr_a1);
                     assign FpgaPins_Fpga_CPU_rs2_valid_a1   = !FpgaPins_Fpga_CPU_reset_a1 & (FpgaPins_Fpga_CPU_is_r_instr_a1 | FpgaPins_Fpga_CPU_is_s_instr_a1 | FpgaPins_Fpga_CPU_is_b_instr_a1);
            
                  //_@2 // Operand Selection
                     assign FpgaPins_Fpga_CPU_rf_rd_en1_a2 = FpgaPins_Fpga_CPU_rs1_valid_a2;
                     assign FpgaPins_Fpga_CPU_rf_rd_en2_a2 = FpgaPins_Fpga_CPU_rs2_valid_a2;
                     assign FpgaPins_Fpga_CPU_rf_rd_index1_a2[4:0] = FpgaPins_Fpga_CPU_rs1_a2;
                     assign FpgaPins_Fpga_CPU_rf_rd_index2_a2[4:0] = FpgaPins_Fpga_CPU_rs2_a2;
            
                     assign FpgaPins_Fpga_CPU_src1_value_a2[31:0] = (FpgaPins_Fpga_CPU_rf_wr_en_a3 && (FpgaPins_Fpga_CPU_rd_a3 == FpgaPins_Fpga_CPU_rs1_a2)) ? FpgaPins_Fpga_CPU_rf_wr_data_a3 : FpgaPins_Fpga_CPU_rf_rd_data1_a2;
                     assign FpgaPins_Fpga_CPU_src2_value_a2[31:0] = (FpgaPins_Fpga_CPU_rf_wr_en_a3 && (FpgaPins_Fpga_CPU_rd_a3 == FpgaPins_Fpga_CPU_rs2_a2)) ? FpgaPins_Fpga_CPU_rf_wr_data_a3 : FpgaPins_Fpga_CPU_rf_rd_data2_a2;
            
                     assign FpgaPins_Fpga_CPU_alu_op1_a2[31:0] =
                        FpgaPins_Fpga_CPU_is_auipc_a2 | FpgaPins_Fpga_CPU_is_jump_a2 ? FpgaPins_Fpga_CPU_pc_a2 :
                                               FpgaPins_Fpga_CPU_src1_value_a2;
                     assign FpgaPins_Fpga_CPU_alu_op2_a2[31:0] =
                        FpgaPins_Fpga_CPU_is_r_instr_a2 || FpgaPins_Fpga_CPU_is_b_instr_a2 ? FpgaPins_Fpga_CPU_src2_value_a2 :
                        FpgaPins_Fpga_CPU_is_jump_a2                   ? 32'h0000_0004 :
                                                     FpgaPins_Fpga_CPU_imm_a2;
            
                     assign FpgaPins_Fpga_CPU_tgt_pc_op1_a2[31:0] = FpgaPins_Fpga_CPU_is_jalr_a2 ? FpgaPins_Fpga_CPU_src1_value_a2 : FpgaPins_Fpga_CPU_pc_a2;
                     assign FpgaPins_Fpga_CPU_tgt_pc_op2_a2[31:0] = FpgaPins_Fpga_CPU_imm_a2;
            
                  //_@3 // Execute, Register Write
                     assign FpgaPins_Fpga_CPU_valid_a3 = !FpgaPins_Fpga_CPU_reset_a3 && !(FpgaPins_Fpga_CPU_valid_taken_br_a4 || FpgaPins_Fpga_CPU_valid_taken_br_a5 || FpgaPins_Fpga_CPU_valid_load_a4 || FpgaPins_Fpga_CPU_valid_load_a5 || FpgaPins_Fpga_CPU_valid_jump_a4 || FpgaPins_Fpga_CPU_valid_jump_a5);
                     assign FpgaPins_Fpga_CPU_valid_load_a3  = FpgaPins_Fpga_CPU_is_load_a3  && FpgaPins_Fpga_CPU_valid_a3;
                     assign FpgaPins_Fpga_CPU_valid_store_a3 = FpgaPins_Fpga_CPU_is_store_a3 && FpgaPins_Fpga_CPU_valid_a3;
                     assign FpgaPins_Fpga_CPU_valid_jump_a3  = FpgaPins_Fpga_CPU_is_jump_a3  && FpgaPins_Fpga_CPU_valid_a3;
                     assign FpgaPins_Fpga_CPU_valid_taken_br_a3 =
                        !FpgaPins_Fpga_CPU_valid_a3  ? 1'b0 :
                        FpgaPins_Fpga_CPU_is_beq_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 == FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_bne_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 != FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_bltu_a3 ? FpgaPins_Fpga_CPU_result_a3[0] :
                        FpgaPins_Fpga_CPU_is_bgeu_a3 ? !FpgaPins_Fpga_CPU_result_a3[0] :
                        FpgaPins_Fpga_CPU_is_blt_a3  ? FpgaPins_Fpga_CPU_result_a3[0] :
                        FpgaPins_Fpga_CPU_is_bge_a3  ? !FpgaPins_Fpga_CPU_result_a3[0] :
                                   1'b0;
                     assign FpgaPins_Fpga_CPU_valid_tgt_pc_a3 = FpgaPins_Fpga_CPU_valid_taken_br_a3 | FpgaPins_Fpga_CPU_valid_jump_a3;
            
                     // Target PC Adder
                     assign FpgaPins_Fpga_CPU_tgt_pc_a3[31:0] = FpgaPins_Fpga_CPU_tgt_pc_op1_a3 + FpgaPins_Fpga_CPU_tgt_pc_op2_a3;
            
                     // ALU
                     assign FpgaPins_Fpga_CPU_sra_result_a3[63:0] = { {32{FpgaPins_Fpga_CPU_alu_op1_a3[31]}}, FpgaPins_Fpga_CPU_alu_op1_a3} >> FpgaPins_Fpga_CPU_alu_op2_a3[4:0];
                     assign FpgaPins_Fpga_CPU_sltu_result_a3[31:0] = FpgaPins_Fpga_CPU_alu_op1_a3 < FpgaPins_Fpga_CPU_alu_op2_a3 ? 32'h0000_0001 : 32'h0000_0000;
                     assign FpgaPins_Fpga_CPU_result_a3[31:0] =
                        FpgaPins_Fpga_CPU_is_add_op_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 + FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_and_op_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 & FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_lui_a3     ? {FpgaPins_Fpga_CPU_alu_op2_a3[31:12], 12'h000} :
                        FpgaPins_Fpga_CPU_is_or_op_a3   ? FpgaPins_Fpga_CPU_alu_op1_a3 | FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_sll_op_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 << FpgaPins_Fpga_CPU_alu_op2_a3[4:0] :
                        FpgaPins_Fpga_CPU_is_slt_op_a3  ? ((FpgaPins_Fpga_CPU_alu_op1_a3[31] == FpgaPins_Fpga_CPU_alu_op2_a3[31]) ? FpgaPins_Fpga_CPU_sltu_result_a3 : (FpgaPins_Fpga_CPU_alu_op1_a3[31] == 1'b1 ? 32'h0000_0001 : 32'h0000_0000)) :
                        FpgaPins_Fpga_CPU_is_sltu_op_a3 ? FpgaPins_Fpga_CPU_sltu_result_a3 :
                        FpgaPins_Fpga_CPU_is_sra_op_a3  ? FpgaPins_Fpga_CPU_sra_result_a3[31:0] :
                        FpgaPins_Fpga_CPU_is_srl_op_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 >> FpgaPins_Fpga_CPU_alu_op2_a3[4:0] :
                        FpgaPins_Fpga_CPU_is_sub_a3     ? FpgaPins_Fpga_CPU_alu_op1_a3 - FpgaPins_Fpga_CPU_alu_op2_a3 :
                        FpgaPins_Fpga_CPU_is_xor_op_a3  ? FpgaPins_Fpga_CPU_alu_op1_a3 ^ FpgaPins_Fpga_CPU_alu_op2_a3 :
                                      32'hxxxx_xxxx;
            
                     // Register Write
                     assign FpgaPins_Fpga_CPU_rf_wr_en_a3 = (FpgaPins_Fpga_CPU_valid_a3 && FpgaPins_Fpga_CPU_rd_valid_a3 && (FpgaPins_Fpga_CPU_rd_a3 != 5'h00) && !FpgaPins_Fpga_CPU_valid_load_a3) || FpgaPins_Fpga_CPU_valid_load_a5;
                     assign FpgaPins_Fpga_CPU_rf_wr_index_a3[4:0] = FpgaPins_Fpga_CPU_valid_a3 ? FpgaPins_Fpga_CPU_rd_a3 : FpgaPins_Fpga_CPU_rd_a5;
                     assign FpgaPins_Fpga_CPU_rf_wr_data_a3[31:0] = FpgaPins_Fpga_CPU_valid_a3 ? FpgaPins_Fpga_CPU_result_a3 : FpgaPins_Fpga_CPU_ld_data_a5;
            
                  //_@4 // Data Memory R/W
                     assign dmem_rd_en = FpgaPins_Fpga_CPU_valid_load_a4;
                     assign dmem_wr_en = FpgaPins_Fpga_CPU_valid_store_a4;
                     assign dmem_addr = FpgaPins_Fpga_CPU_result_a4[DMEM_BYTE_ADDR_WIDTH-1:2];
                     assign dmem_wr_byte_en = 4'b1111; // Just implement LW/SW for now
                     assign dmem_wr_data = FpgaPins_Fpga_CPU_src2_value_a4;
                     assign FpgaPins_Fpga_CPU_ld_data_a4[31:0] = dmem_rd_data;
            
                  // Note that pipesignals assigned here can be found under /fpga_pins/fpga.
            
            
            
            
               // Assert these to end simulation (before Makerchip cycle limit).
               // Note, for Makerchip simulation these are passed in uo_out to top-level module's passed/failed signals.
               //*passed = *top.cyc_cnt > 40;
               //*passed = (|cpu/xreg[15]>>5$value == (1+2+3+4+5+6+7+8+9)) && (*top.cyc_cnt > 65);
               //*passed = |cpu/xreg[15]>>5$value == (1+2+3+4+5+6+7+8+9);
               //*failed = 1'b0;
            
               // Connect Tiny Tapeout outputs. Note that uio_ outputs are not available in the Tiny-Tapeout-3-based FPGA boards.
               // *uo_out = {6'b0, *failed, *passed};
               // assign uio_out = 8'b0;
               // assign uio_oe = 8'b0;
            
               // Macro instantiations to be uncommented when instructed for:
               //  o instruction memory
               //  o register file
               //  o data memory
               //  o CPU visualization
               //_|cpu
                  // m4+imem(@1)    // Args: (read stage)
                  //_\source /raw.githubusercontent.com/efabless/chipcraftmestcourse/main/tlvlib/riscvshelllib.tlv 33   // Instantiated from top.tlv, 291 as: m4+rf(@2, @3)
                     // Reg File
                     //_@3
                        for (xreg = 0; xreg <= 15; xreg++) begin : L1_FpgaPins_Fpga_CPU_Xreg //_/xreg

                           // For $wr.
                           logic L1_wr_a3;

                           assign L1_wr_a3 = FpgaPins_Fpga_CPU_rf_wr_en_a3 && (FpgaPins_Fpga_CPU_rf_wr_index_a3 != 5'b0) && (FpgaPins_Fpga_CPU_rf_wr_index_a3 == xreg);
                           assign FpgaPins_Fpga_CPU_Xreg_value_a3[xreg][31:0] = FpgaPins_Fpga_CPU_reset_a3 ?   xreg           :
                                          L1_wr_a3        ?   FpgaPins_Fpga_CPU_rf_wr_data_a3 :
                                                         FpgaPins_Fpga_CPU_Xreg_value_a4[xreg][31:0];
                        end
                     //_@2
                        //_?$rf_rd_en1
                           assign FpgaPins_Fpga_CPU_rf_rd_data1_a2[31:0] = FpgaPins_Fpga_CPU_Xreg_value_a4[FpgaPins_Fpga_CPU_rf_rd_index1_a2[3:0]];
                        //_?$rf_rd_en2
                           assign FpgaPins_Fpga_CPU_rf_rd_data2_a2[31:0] = FpgaPins_Fpga_CPU_Xreg_value_a4[FpgaPins_Fpga_CPU_rf_rd_index2_a2[3:0]];
                        `BOGUS_USE(FpgaPins_Fpga_CPU_rf_rd_data1_a2 FpgaPins_Fpga_CPU_rf_rd_data2_a2)
                  //_\end_source  // Args: (read stage, write stage) - if equal, no register bypass is required
                  // m4+dmem(@4)    // Args: (read/write stage)
            
               // m4+cpu_viz(@4)    // For visualisation, argument should be at least equal to the last stage of CPU logic. @4 would work for all labs.
            //_\end_source
   
      // LEDs.
      
   
      // 7-Segment
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 395   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 346 as: m4+fpga_sseg.
         for (digit = 0; digit <= 0; digit++) begin : L1_Digit //_/digit
            
            for (leds = 0; leds <= 7; leds++) begin : L2_Leds //_/leds

               // For $viz_lit.
               logic L2_viz_lit_a0;

               assign L2_viz_lit_a0 = (! L0_sseg_digit_n_a0[digit]) && ! ((leds == 7) ? L0_sseg_decimal_point_n_a0 : L0_sseg_segment_n_a0[leds % 7]);
               
            end
         end
      //_\end_source
   
      // slideswitches
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 454   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 349 as: m4+fpga_switch.
         for (switch = 0; switch <= 7; switch++) begin : L1_Switch //_/switch

            // For $viz_switch.
            logic L1_viz_switch_a0;

            assign L1_viz_switch_a0 = L0_slideswitch_a0[switch];
            
         end
      //_\end_source
   
      // pushbuttons
      
   //_\end_source
   // Label the switch inputs [0..7] (1..8 on the physical switch panel) (top-to-bottom).
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/35e36bd144fddd75495d4cbc01c4fc50ac5bde6f/tlvlib/tinytapeoutlib.tlv 82   // Instantiated from top.tlv, 405 as: m5+tt_input_labels_viz(⌈"UNUSED", "UNUSED", "UNUSED", "UNUSED", "UNUSED", "UNUSED", "UNUSED", "UNUSED"⌉)
      for (input_label = 0; input_label <= 7; input_label++) begin : L1_InputLabel //_/input_label
         
      end
   //_\end_source

//_\SV
endmodule


// Undefine macros defined by SandPiper.
`undef BOGUS_USE

module synchronizer (
   input  logic clk,    //your local clock
   input  logic async,  //unsynchronized signal
   output logic sync); //synchronized signal

   // Create a signal buffer
   logic [1:0] buff;

   always_ff @ (posedge clk) 
      buff <= {buff[0], async};

   assign sync = buff[1];

endmodule

module neg_edge_detector (
   input  logic clk,
   input  logic rst,
   input  logic signal_in,
   output logic edge_detected);

   logic register;

   always_ff @(posedge clk) begin
      if (rst) register <= 1;
      else register <= signal_in;
   end

   assign edge_detected = register & ~signal_in;

endmodule

module pos_edge_detector (
   input  logic clk,
   input  logic rst,
   input  logic signal_in,
   output logic edge_detected);

   logic register;

   always_ff @(posedge clk) begin
      if (rst) register <= 1;
      else register <= signal_in;
   end

   assign edge_detected = ~register & signal_in;

endmodule

module shift_register #(
   parameter int unsigned NUM_BITS = 8,
   parameter int unsigned RST_VALUE = 0)
(
   input  logic clk,
   input  logic rst,
   input  logic serial_in,
   input  logic shift_enable,
   input  logic [NUM_BITS-1:0] parallel_in,
   input  logic load_enable,
   output logic serial_out,
   output logic [NUM_BITS-1:0] parallel_out);

   logic [NUM_BITS-1:0] register;

   always_ff @(posedge clk) begin
      if (rst) register <= RST_VALUE[NUM_BITS-1:0];
      else if (load_enable) register <= parallel_in;
      else if (shift_enable) begin
         for (int unsigned i = 0; i < NUM_BITS-1; i++) register[i] <= register[i+1];
         register[NUM_BITS-1] <= serial_in;
      end
      else register <= register;
   end

   always_comb begin
      parallel_out = register;
      serial_out = register[0];
   end

endmodule

module uart_rx #(
   parameter int unsigned COUNTER_WIDTH = 24)
(
   input  logic clk,
   input  logic rst,
   input  logic uart_rx_in,
   output logic [7:0] data,                         // Valid only when "ready" is high, undefined otherwise
   output logic [COUNTER_WIDTH-1:0] cycles_per_bit, // Length of the first packet starting bit in clock cycles
   output ready);                                   // Held high for duration of STOP bit, low all other times

   // Declare intermediate wires
   logic baud_rate_known, uart_rx_in_synced, start_detected, rising_edge, timer_rst, half_bit, full_bit, shift_en;
   logic [COUNTER_WIDTH-1:0] counter_val;
   enum logic [3:0] {
      STATE_IDLE  = 4'h0,
      STATE_START = 4'h1,
      STATE_D0    = 4'h2,
      STATE_D1    = 4'h3,
      STATE_D2    = 4'h4,
      STATE_D3    = 4'h5,
      STATE_D4    = 4'h6,
      STATE_D5    = 4'h7,
      STATE_D6    = 4'h8,
      STATE_D7    = 4'h9,
      STATE_STOP  = 4'hA
   } state;

   // Upon Reset, Baud Rate is not known
   always_ff @(posedge clk) begin
      if (rst) baud_rate_known <= 1'b0;
      else if ((state == STATE_STOP) && (start_detected || full_bit)) baud_rate_known <= 1'b1;
   end

   // Connect synchronizer
   synchronizer uart_rx_in_synchronizer(
      .clk(clk),
      .async(uart_rx_in),
      .sync(uart_rx_in_synced));

   // Connect edge detectors
   neg_edge_detector start_detector(
      .clk(clk),
      .rst(rst),
      .signal_in(uart_rx_in_synced),
      .edge_detected(start_detected));
   pos_edge_detector rising_edge_detector(
      .clk(clk),
      .rst(rst),
      .signal_in(uart_rx_in_synced),
      .edge_detected(rising_edge));

   // Connect shift register
   assign shift_en = ((state > STATE_START) && (state < STATE_STOP) && half_bit && baud_rate_known) ? 1'b1:1'b0;
   shift_register #(
      .NUM_BITS(8),
      .RST_VALUE(0))
   shift_reg(
      .clk(clk),
      .rst(rst),
      .serial_in(uart_rx_in_synced),
      .shift_enable(shift_en),
      .parallel_in(8'h0),
      .load_enable(1'b0),
      .serial_out(),
      .parallel_out(data));

   // Implement timer
   assign timer_rst = ((state == STATE_IDLE) || (state == STATE_STOP && start_detected) || full_bit || rst) ? 1'b1:1'b0;
   assign half_bit = counter_val == cycles_per_bit >> 1 ? 1'b1 : 1'b0;
   assign full_bit = (counter_val >= cycles_per_bit) || (state == STATE_START && !baud_rate_known && rising_edge) ? 1'b1 : 1'b0;
   always_ff @(posedge clk) begin
      if (rst) cycles_per_bit <= {COUNTER_WIDTH{1'b1}};
      else if (state == STATE_START && rising_edge) cycles_per_bit <= counter_val;
   end
   always_ff @(posedge clk) begin
      if (timer_rst) counter_val <= '0;
      else counter_val <= counter_val + 1;
   end

   // State machine logic
   always_ff @(posedge clk) begin
      if (rst || (state > STATE_STOP)) state <= STATE_IDLE;
      else if (start_detected && (state == STATE_IDLE || state == STATE_STOP)) state <= STATE_START;
      else if (full_bit)
         case (state)
            STATE_START:    state <= STATE_D0;
            STATE_D0:       state <= STATE_D1;
            STATE_D1:       state <= STATE_D2;
            STATE_D2:       state <= STATE_D3;
            STATE_D3:       state <= STATE_D4;
            STATE_D4:       state <= STATE_D5;
            STATE_D5:       state <= STATE_D6;
            STATE_D6:       state <= STATE_D7;
            STATE_D7:       state <= STATE_STOP;
            STATE_STOP:     state <= STATE_IDLE;
            default:        state <= state;
         endcase
      else state <= state;
   end

   // Connect outputs
   assign ready = (state == STATE_STOP && baud_rate_known) ? 1'b1:1'b0;

endmodule

module uart_tx #(
   parameter int unsigned COUNTER_WIDTH = 24)
(
   input  logic clk,
   input  logic rst,
   output logic uart_tx_out,
   input  logic [7:0] data,
   input  logic req,
   input  logic [COUNTER_WIDTH-1:0] cycles_per_bit,
   output logic empty,
   output logic error);

   // Declare intermediate wires
   logic full_bit, idle_state;
   logic [COUNTER_WIDTH-1:0] counter_val;
   enum logic [3:0] {
      STATE_IDLE  = 4'h0,
      STATE_START = 4'h1,
      STATE_D0    = 4'h2,
      STATE_D1    = 4'h3,
      STATE_D2    = 4'h4,
      STATE_D3    = 4'h5,
      STATE_D4    = 4'h6,
      STATE_D5    = 4'h7,
      STATE_D6    = 4'h8,
      STATE_D7    = 4'h9,
      STATE_STOP  = 4'hA
   } state;

   assign idle_state = (state == STATE_IDLE) ? 1'b1:1'b0;

   // Connect shift register
   shift_register #(
      .NUM_BITS(9),
      .RST_VALUE(1))
   shift_reg(
      .clk(clk),
      .rst(rst),
      .serial_in(1'b1),
      .shift_enable(full_bit),
      .parallel_in({data, 1'b0}),
      .load_enable(idle_state & req),
      .serial_out(uart_tx_out),
      .parallel_out());

   // Implement timer
   assign full_bit = (counter_val >= cycles_per_bit) ? 1'b1 : 1'b0;
   always_ff @(posedge clk) begin
      if (full_bit || idle_state || rst) counter_val <= '0;
      else counter_val <= counter_val + 1;
   end

   // State machine logic
   always_ff @(posedge clk) begin
      if (rst || (state > STATE_STOP)) state <= STATE_IDLE;
      else if (idle_state & req) state <= STATE_START;
      else if (full_bit)
         case (state)
            STATE_START:    state <= STATE_D0;
            STATE_D0:       state <= STATE_D1;
            STATE_D1:       state <= STATE_D2;
            STATE_D2:       state <= STATE_D3;
            STATE_D3:       state <= STATE_D4;
            STATE_D4:       state <= STATE_D5;
            STATE_D5:       state <= STATE_D6;
            STATE_D6:       state <= STATE_D7;
            STATE_D7:       state <= STATE_STOP;
            STATE_STOP:     state <= STATE_IDLE;
            default:        state <= STATE_IDLE;
         endcase
      else state <= state;
   end

   // Connect outputs
   assign empty = idle_state;
   assign error = ~idle_state & req;

endmodule

module uart_ctrl #(
   parameter int unsigned IMEM_BYTE_ADDR_WIDTH = 6, // 64 bytes of storage, or 16 four-byte words
   parameter int unsigned DMEM_BYTE_ADDR_WIDTH = 6) // 64 bytes of storage, or 16 four-byte words
(
   input  logic clk,
   input  logic rst,
   input  logic rx_ready,
   input  logic tx_empty,
   input  logic tx_error,
   output logic cpu_rst,
   output logic tx_req,
   output logic imem_ctrl,
   output logic imem_wr_en,
   output logic [IMEM_BYTE_ADDR_WIDTH-1:0] imem_addr,
   output logic dmem_ctrl,
   output logic dmem_rd_en,
   output logic [DMEM_BYTE_ADDR_WIDTH-1:0] dmem_addr);

   localparam int unsigned NUM_IMEM_BYTES = 2**IMEM_BYTE_ADDR_WIDTH;
   localparam int unsigned NUM_DMEM_BYTES = 2**DMEM_BYTE_ADDR_WIDTH;

   // Declare intermediate wires
   logic rd_complete, wr_data_ready, all_imem_written;
   enum logic [1:0] {
      STATE_RESET      = 2'b00,
      STATE_DATA_WRITE = 2'b01,
      STATE_IDLE       = 2'b10,
      STATE_DATA_READ  = 2'b11
   } state;

   // Assign intermediate wires
   /* verilator lint_off WIDTHEXPAND */
   assign rd_complete = ((state == STATE_DATA_READ) && (dmem_addr == NUM_DMEM_BYTES-1) && dmem_rd_en) ? 1'b1 : 1'b0;
   assign all_imem_written = ((state == STATE_DATA_WRITE) && (imem_addr == NUM_IMEM_BYTES-1) && imem_wr_en) ? 1'b1 : 1'b0;
   /* verilator lint_on WIDTHEXPAND */
   pos_edge_detector wr_data_ready_detect (
      .clk(clk),
      .rst(rst),
      .signal_in(rx_ready),
      .edge_detected(wr_data_ready)
   );

   // State machine logic
   always_ff @(posedge clk) begin
      if (rst) state <= STATE_RESET;
      else begin
         case (state)
            STATE_RESET:      if (!rst)             state <= STATE_DATA_WRITE;
            STATE_DATA_WRITE: if (all_imem_written) state <= STATE_IDLE;
            STATE_IDLE:       if (wr_data_ready)    state <= STATE_DATA_READ;
            STATE_DATA_READ:  if (rd_complete)      state <= STATE_IDLE;
         endcase
      end // else
   end // always_ff

   // I-Memory Address Counter
   always_ff @(posedge clk) begin
      if (rst) imem_addr <= '0;
      else if (state == STATE_RESET) imem_addr <= '0;
      else if (state == STATE_IDLE)  imem_addr <= '0;
      else if (state == STATE_DATA_WRITE && imem_wr_en) imem_addr <= imem_addr + 1;
   end //always_ff

   // D-Memory Address Counter
   always_ff @(posedge clk) begin
      if (rst) dmem_addr <= '0;
      else if (state == STATE_RESET) dmem_addr <= '0;
      else if (state == STATE_IDLE)  dmem_addr <= '0;
      else if (state == STATE_DATA_READ && dmem_rd_en) dmem_addr <= dmem_addr + 1;
   end //always_ff

   // Connect outputs
   assign cpu_rst    = (state == STATE_RESET || state == STATE_DATA_WRITE || rst) ? 1'b1 : 1'b0;
   assign imem_ctrl  = cpu_rst;
   assign dmem_ctrl  = cpu_rst;
   assign dmem_rd_en = (state == STATE_DATA_READ && tx_empty) ? 1'b1 : 1'b0;
   assign imem_wr_en = (state == STATE_DATA_WRITE && wr_data_ready) ? 1'b1 : 1'b0;
   assign tx_req     = dmem_rd_en;

endmodule

module mem_rf #(
   parameter int unsigned MEM_BYTE_ADDR_WIDTH = 6) // 64 bytes of storage, or 16 four-byte words
(
   input  logic clk,
   input  logic rst,
   // UART Memory Interface
   input  logic umem_ctrl,
   input  logic umem_rd_en,
   input  logic umem_wr_en,
   input  logic [MEM_BYTE_ADDR_WIDTH-1:0] umem_addr,
   input  logic [7:0] umem_wr_data,
   output logic [7:0] umem_rd_data,
   // CPU Memory Interface
   input  logic cpu_mem_rd_en,
   input  logic cpu_mem_wr_en,
   input  logic [MEM_BYTE_ADDR_WIDTH-3:0] cpu_mem_addr, // Two fewer bits than umem since addressing 4 byte values
   input  logic [3:0] cpu_mem_wr_byte_en,
   input  logic [31:0] cpu_mem_wr_data,
   output logic [31:0] cpu_mem_rd_data);

   localparam int unsigned NUM_MEM_BYTES = 2**MEM_BYTE_ADDR_WIDTH;

   logic [7:0] reg_file [NUM_MEM_BYTES];

   always_ff @(posedge clk) begin
      if (rst) begin
         for (int unsigned i = 0; i < NUM_MEM_BYTES; i++) reg_file[i] = 8'h00;
      end // if
      else if (umem_ctrl && umem_wr_en)
         reg_file[umem_addr] <= umem_wr_data;
      else if (!umem_ctrl && cpu_mem_wr_en) begin
         if (cpu_mem_wr_byte_en[3]) reg_file[{cpu_mem_addr, 2'b11}] <= cpu_mem_wr_data[31:24];
         if (cpu_mem_wr_byte_en[2]) reg_file[{cpu_mem_addr, 2'b10}] <= cpu_mem_wr_data[23:16];
         if (cpu_mem_wr_byte_en[1]) reg_file[{cpu_mem_addr, 2'b01}] <= cpu_mem_wr_data[15:8];
         if (cpu_mem_wr_byte_en[0]) reg_file[{cpu_mem_addr, 2'b00}] <= cpu_mem_wr_data[7:0];
      end
   end // always_ff

   assign umem_rd_data = reg_file[umem_addr];
   assign cpu_mem_rd_data =
      {reg_file[{cpu_mem_addr, 2'b11}],
       reg_file[{cpu_mem_addr, 2'b10}],
       reg_file[{cpu_mem_addr, 2'b01}],
       reg_file[{cpu_mem_addr, 2'b00}]};

endmodule

module uart_top #(
   parameter int unsigned COUNTER_WIDTH = 24,
   parameter int unsigned IMEM_BYTE_ADDR_WIDTH = 6, // 64 bytes of storage, or 16 four-byte words
   parameter int unsigned DMEM_BYTE_ADDR_WIDTH = 6) // 64 bytes of storage, or 16 four-byte words
(
   input  logic clk,
   // User Interface
   input  logic rst,
   input  logic rx_in,
   output logic tx_out,
   // CPU Interface
   output logic cpu_rst,
   input  logic imem_rd_en,
   input  logic [IMEM_BYTE_ADDR_WIDTH-3:0] imem_rd_addr,
   output logic [31:0] imem_rd_data,
   input  logic dmem_rd_en,
   input  logic dmem_wr_en,
   input  logic [DMEM_BYTE_ADDR_WIDTH-3:0] dmem_addr,
   input  logic [3:0] dmem_wr_byte_en,
   input  logic [31:0] dmem_wr_data,
   output logic [31:0] dmem_rd_data);

   logic rx_ready, tx_empty, tx_error, tx_req, imem_uart_ctrl, imem_uart_wr_en, dmem_uart_ctrl, dmem_uart_rd_en;
   logic [IMEM_BYTE_ADDR_WIDTH-1:0] imem_uart_addr;
   logic [DMEM_BYTE_ADDR_WIDTH-1:0] dmem_uart_addr;
   logic [7:0] umem_rd_data, umem_wr_data;
   logic [COUNTER_WIDTH-1:0] cycles_per_bit;

   uart_rx #(
      .COUNTER_WIDTH(COUNTER_WIDTH))
   uart_rx0 (
      .clk(clk),
      .rst(rst),
      .uart_rx_in(rx_in),
      .data(umem_wr_data),
      .cycles_per_bit(cycles_per_bit),
      .ready(rx_ready));

   uart_tx #(
      .COUNTER_WIDTH(COUNTER_WIDTH))
   uart_tx0 (
      .clk(clk),
      .rst(rst),
      .uart_tx_out(tx_out),
      .data(umem_rd_data),
      .req(tx_req),
      .cycles_per_bit(cycles_per_bit),
      .empty(tx_empty),
      .error(tx_error));

   uart_ctrl #(
      .IMEM_BYTE_ADDR_WIDTH(IMEM_BYTE_ADDR_WIDTH),
      .DMEM_BYTE_ADDR_WIDTH(DMEM_BYTE_ADDR_WIDTH))
   uart_ctrl0 (
      .clk(clk),
      .rst(rst),
      .rx_ready(rx_ready),
      .tx_empty(tx_empty),
      .tx_error(tx_error),
      .cpu_rst(cpu_rst),
      .tx_req(tx_req),
      .imem_ctrl(imem_uart_ctrl),
      .imem_wr_en(imem_uart_wr_en),
      .imem_addr(imem_uart_addr),
      .dmem_ctrl(dmem_uart_ctrl),
      .dmem_rd_en(dmem_uart_rd_en),
      .dmem_addr(dmem_uart_addr));

   mem_rf #(
      .MEM_BYTE_ADDR_WIDTH(IMEM_BYTE_ADDR_WIDTH))
   imem0 (
      .clk(clk),
      .rst(rst),
      .umem_ctrl(imem_uart_ctrl),
      .umem_rd_en(0),
      .umem_wr_en(imem_uart_wr_en),
      .umem_addr(imem_uart_addr),
      .umem_wr_data(umem_wr_data),
      .umem_rd_data(),
      .cpu_mem_rd_en(imem_rd_en),
      .cpu_mem_wr_en(0),
      .cpu_mem_addr(imem_rd_addr),
      .cpu_mem_wr_byte_en('0),
      .cpu_mem_wr_data('0),
      .cpu_mem_rd_data(imem_rd_data));

   mem_rf #(
      .MEM_BYTE_ADDR_WIDTH(DMEM_BYTE_ADDR_WIDTH))
   dmem0 (
      .clk(clk),
      .rst(rst),
      .umem_ctrl(dmem_uart_ctrl),
      .umem_rd_en(dmem_uart_rd_en),
      .umem_wr_en(0),
      .umem_addr(dmem_uart_addr),
      .umem_wr_data('0),
      .umem_rd_data(umem_rd_data),
      .cpu_mem_rd_en(dmem_rd_en),
      .cpu_mem_wr_en(dmem_wr_en),
      .cpu_mem_addr(dmem_addr),
      .cpu_mem_wr_byte_en(dmem_wr_byte_en),
      .cpu_mem_wr_data(dmem_wr_data),
      .cpu_mem_rd_data(dmem_rd_data));
endmodule
